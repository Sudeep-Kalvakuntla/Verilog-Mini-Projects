module uut(
  reg A0,
  reg A1,
  reg A2,
  reg A3,
  wire Y
);

endmodule
